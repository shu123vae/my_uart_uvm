`ifndef MY_TRANSACTION
`define MY_TRANSACTION

`include "uvm_macros.svh"
import uvm_pkg::*;

class my_transaction extends uvm_sequence_item;

	bit [7:0] SerDataIn=8'h5A;	//in
	rand bit SerInParity;		//in
	rand bit inject_error;	//in
	bit [8:0] PalDataOut;	//out
	bit PalDataOutValid;	//out


	bit [7:0] PalDataIn=8'hA1;//in
	bit PalDataInEn;	//in
	bit PalDataInPermit;	//out
	bit [7:0] SerDataOut;	//out


constraint c_parity{
    SerInParity == ~^SerDataIn;
    if (inject_error) 
	SerInParity != ~^SerDataIn;
}

`uvm_object_utils_begin(my_transaction)
	`uvm_field_int(SerDataIn,UVM_ALL_ON)
	`uvm_field_int(PalDataOut,UVM_ALL_ON)
	`uvm_field_int(PalDataOutValid,UVM_ALL_ON)
	`uvm_field_int(PalDataIn, UVM_ALL_ON)
	`uvm_field_int(PalDataInEn, UVM_ALL_ON)	
	`uvm_field_int(PalDataInPermit, UVM_ALL_ON)
	`uvm_field_int(SerDataOut, UVM_ALL_ON)
`uvm_object_utils_end

function new(string name="my_transaction");
	super.new(name);
	`uvm_info("my_transaction","the my_transaction new is called!",UVM_LOW)
endfunction

endclass

`endif